`timescale 1ns/1ns

module mvs_cart(
	input nRESET,
	input CLK_24M, CLK_12M, CLK_8M, CLK_68KCLKB, CLK_4MB,
	
	input nAS, M68K_RW,
	input [19:1] M68K_ADDR,
	inout [15:0] M68K_DATA,
	input nROMOE, nROMOEL, nROMOEU,
	input nPORTADRS, nPORTOEL, nPORTOEU, nPORTWEL, nPORTWEU, 
	output nROMWAIT, nPWAIT0, nPWAIT1, PDTACK,
	
	input nSLOTCS,
	
	input [23:0] PBUS,
	input CA4,
	input S2H1,
	input PCK1B,
	input PCK2B,
	output [31:0] CR,
	output [7:0] FIXD,
	
	inout [7:0] SDRAD,
	input [9:8] SDRA_L,
	input [23:20] SDRA_U,
	input SDRMPX, nSDROE,
	
	inout [7:0] SDPAD,
	input [11:8] SDPA,
	input SDPMPX, nSDPOE,
	
	input SDRD0, SDRD1, nSDROM, nSDMRD,
	input [15:0] SDA,
	inout [7:0] SDD
);
	
	prog_board PROG(nSDROE, SDRMPX, SDRA_U, SDRA_L, nSDPOE, SDPMPX, SDPA, nSLOTCS, nPORTADRS, nPORTWEL, nPORTWEU,
						nPORTOEL, nPORTOEU, nROMOEL, nROMOEU, nAS, M68K_RW, M68K_DATA, M68K_ADDR, CLK_68KCLKB, nROMWAIT,
						nPWAIT0, nPWAIT1, PDTACK, nROMOE, CLK_4MB, nRESET, SDPAD, SDRAD);
	
	cha_board CHA(SDA, nSLOTCS, CR, CA4, S2H1, PCK2B, PCK1B, PBUS, CLK_24M, CLK_12M, CLK_8M, nRESET, FIXD,
						SDRD0, SDRD1, nSDROM, nSDMRD, SDD);

endmodule
