`timescale 1ns/1ns

module ym_fm(
	input PHI_S
);

	always @(posedge PHI_S)		// posedge ?
	begin
		// Todo...
	end
	
endmodule
