// NeoGeo logic definition (simulation only)
// Copyright (C) 2018 Sean Gonsalves
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.

`timescale 1ns/1ns

module resetp(
	input CLK_24MB,
	input RESET,
	output RESETP
);

	// nRESET  ""|_________|""""""
	// nRESETP """"""""""""""|_|""
	
	FDM O52(CLK_24MB, RESET, O52_Q, );
	FDM O49(CLK_24MB, O52_Q, , O49_nQ);
	
	assign RESETP = ~&{O49_nQ, O52_Q};
	
endmodule
